`timescale 1ns / 1ps
`include "uvm_macros.svh"
import uvm_pkg::*;

class apb_config extends uvm_object;
	`uvm_object_utils(apb_config)

	function new(string path = "apb_config");
		super.new(path);
	endfunction

	uvm_active_passive_enum is_active = UVM_ACTIVE;

endclass

typedef enum bit[1:0] {readd = 0, writed = 1, rst = 2} oper_mode;

class transaction extends uvm_sequence_item;

	rand oper_mode op;

  	randc logic [31:0] paddr;
  	rand logic pwrite;
  	rand logic [31:0] pwdata;


	logic [31:0] prdata;
  	logic pslverr;
  	logic pready;

	function new(input string path = "transaction");
		super.new(path);
	endfunction

	`uvm_object_utils_begin(transaction)

	`uvm_field_int(paddr,UVM_DEFAULT)
	`uvm_field_int(pwrite,UVM_DEFAULT)
	`uvm_field_int(pwdata,UVM_DEFAULT)
	`uvm_field_int(prdata,UVM_DEFAULT)
	`uvm_field_int(pslverr,UVM_DEFAULT)
	`uvm_field_int(pready,UVM_DEFAULT)
	`uvm_field_enum(oper_mode, op, UVM_DEFAULT)

	`uvm_object_utils_end

	constraint addr_c {paddr < 32; }
	constraint addr_c_err { paddr >= 32; }

endclass

// write data sequence 
class write_data extends uvm_sequence #(transaction);
	`uvm_object_utils(write_data)

	transaction tr;
	integer i = 15;

	function new(input string path = "write_data");
		super.new(path);
	endfunction


	virtual task body();
		repeat(i) begin

			tr = transaction::type_id::create("tr");
			tr.addr_c.constraint_mode(1);
			tr.addr_c_err.constraint_mode(0);

			start_item(tr);
			assert(tr.randomize()) else 
				`uvm_error("SEQ","Randomization Failed")
			tr.op = writed;
			`uvm_info("SEQ","Data Write Request Sent:",UVM_NONE)
			finish_item(tr);

		end
	endtask
endclass

// write error sequence
class write_err extends uvm_sequence #(transaction);
	`uvm_object_utils(write_err)

	transaction tr;
	integer i = 5;

	function new(input string path = "write_err");
		super.new(path);
	endfunction


	virtual task body();
		repeat(i)
		begin
			tr = transaction::type_id::create("tr");
			tr.addr_c.constraint_mode(0);
			tr.addr_c_err.constraint_mode(1);

			start_item(tr);
			assert(tr.randomize())
			else
				`uvm_error("SEQ","Randomization Failed")
			tr.op = writed;
			`uvm_info("SEQ","Illegal Address Data Write Request Sent:",UVM_NONE)
			finish_item(tr);
		end	
	endtask
endclass

//Read Sequence
class read_data extends uvm_sequence #(transaction);
	`uvm_object_utils(read_data)

	transaction tr;
	integer i = 15;

	function new(input string path = "read_data");
		super.new(path);
	endfunction


	virtual task body();
		repeat(i)
		begin
			tr = transaction::type_id::create("tr");
			tr.addr_c.constraint_mode(1);
			tr.addr_c_err.constraint_mode(0);

			start_item(tr);
			assert(tr.randomize())
			else
				`uvm_error("SEQ","Randomization Failed")
			tr.op = readd;
			`uvm_info("SEQ","Data Read Request Sent:",UVM_NONE)
			finish_item(tr);
		end	
	endtask
endclass


//Read Error Sequence
class read_err extends uvm_sequence #(transaction);
	`uvm_object_utils(read_err)

	transaction tr;
	integer i = 5;

	function new(input string path = "read_err");
		super.new(path);
	endfunction


	virtual task body();
		repeat(i)
		begin
			tr = transaction::type_id::create("tr");
			tr.addr_c.constraint_mode(0);
			tr.addr_c_err.constraint_mode(1);

			start_item(tr);
			assert(tr.randomize())
			else
				`uvm_error("SEQ","Randomization Failed")
			tr.op = readd;
			`uvm_info("SEQ","Illegal Address Data Read Request Sent:",UVM_NONE)
			finish_item(tr);
		end	
	endtask
endclass


//Reset Sequence
class reset_dut extends uvm_sequence #(transaction);
	`uvm_object_utils(reset_dut)

	transaction tr;
	integer i = 5;

	function new(input string path = "reset_dut");
		super.new(path);
	endfunction


	virtual task body();
		repeat(i)
		begin
			tr = transaction::type_id::create("tr");
			tr.addr_c.constraint_mode(1);
			tr.addr_c_err.constraint_mode(0);

			start_item(tr);
			assert(tr.randomize())
			else
				`uvm_error("SEQ","Randomization Failed")
			tr.op = rst;
			`uvm_info("SEQ","Reset Request Sent:",UVM_NONE)
			finish_item(tr);
		end	
	endtask
endclass

//Write after read Sequence
class write_read extends uvm_sequence #(transaction);
	`uvm_object_utils(write_read)

	transaction tr;
	integer i = 15;

	function new(input string path = "write_read");
		super.new(path);
	endfunction


	virtual task body();
		repeat(i)
		begin
			tr = transaction::type_id::create("tr");
			tr.addr_c.constraint_mode(1);
			tr.addr_c_err.constraint_mode(0);

			start_item(tr);
			assert(tr.randomize())
			else
				`uvm_error("SEQ","Randomization Failed")
			tr.op = writed;
			`uvm_info("SEQ","Data Write Request Sent:",UVM_NONE)
			finish_item(tr);

			start_item(tr);
			assert(tr.randomize())
			else
				`uvm_error("SEQ","Randomization Failed")
			tr.op = readd;
			`uvm_info("SEQ","Data Read Request Sent:",UVM_NONE)
			finish_item(tr);
		end	
	endtask
endclass



//Read Write bulk Sequence
class writeb_readb extends uvm_sequence #(transaction);
	`uvm_object_utils(writeb_readb)

	transaction tr;
	integer i = 32;

	function new(input string path = "writeb_readb");
		super.new(path);
	endfunction


	virtual task body();
		tr = transaction::type_id::create("tr");
		tr.addr_c.constraint_mode(1);
		tr.addr_c_err.constraint_mode(0);
		repeat(i)
		begin
			start_item(tr);
			assert(tr.randomize())
			else
				`uvm_error("SEQ","Randomization Failed")
			tr.op = writed;
			`uvm_info("SEQ","Data Write Request Sent:",UVM_NONE)
			finish_item(tr);
		end

		tr = transaction::type_id::create("tr");
		tr.addr_c.constraint_mode(1);
		tr.addr_c_err.constraint_mode(0);
		repeat(i)
		begin
			start_item(tr);
			assert(tr.randomize())
			else
				`uvm_error("SEQ","Randomization Failed")
			tr.op = readd;
			`uvm_info("SEQ","Data Read Request Sent:",UVM_NONE)
			finish_item(tr);
		end
	endtask

endclass



class driver extends uvm_driver#(transaction);
	`uvm_component_utils(driver)

	function new(input string path = "driver", input uvm_component parent);
		super.new(path,parent);
	endfunction

	transaction tr;
	virtual apb_if vif;

	virtual function void build_phase(uvm_phase phase);
		super.build_phase(phase);

		tr = transaction::type_id::create("tr");

		if(!uvm_config_db#(virtual apb_if)::get(this,"","vif",vif))
			`uvm_error("DRV","Unable to access Virtual Interface");

	endfunction

	task reset_dut();
		vif.presetn <= 1'b0;
		vif.penable <= 0;
		vif.psel <= 0;
		vif.pwrite <= 0;
		vif.paddr <= 'h0;
		vif.pwdata <= 'h0;
		repeat(5)@(posedge vif.pclk);
		`uvm_info("DRV","Reset Done: Start of Simulation",UVM_NONE);
	endtask

	virtual task run_phase(uvm_phase phase);

		reset_dut();
		forever begin
			seq_item_port.get_next_item(tr);
			
			if(tr.op == rst)
			begin
				vif.presetn <= 1'b0;
				vif.penable <= 0;
				vif.psel <= 0;
				vif.pwrite <= 0;
				vif.paddr <= 'h0;
				vif.pwdata <= 'h0;
				`uvm_info("DRV","Reset done",UVM_NONE);
				@(posedge vif.pclk);

			end

			else if(tr.op == writed)
			begin
				vif.presetn <= 1'b1;
				vif.psel <= 1;
				vif.pwrite <= 1;
				vif.paddr <= tr.paddr;
				vif.pwdata <= tr.pwdata;
				@(posedge vif.pclk);
				vif.penable <= 1;
				@(posedge vif.pready)
				vif.penable <= 0;
				vif.psel <= 0;
				`uvm_info("DRV",$sformatf("Data Write applied to the Interface: Addr = %0d, Wdata = %0d",tr.paddr,tr.pwdata),UVM_NONE);
				@(negedge vif.pready);

			end

			else if(tr.op == readd)
			begin
				vif.presetn <= 1'b1;
				vif.psel <= 1;
				vif.pwrite <= 0;
				vif.paddr <= tr.paddr;
				@(posedge vif.pclk);
				vif.penable <= 1;
				@(posedge vif.pready)
				vif.penable <= 0;
				vif.psel <= 0;
				`uvm_info("DRV",$sformatf("Data Read applied to the Interface: Addr = %0d",tr.paddr),UVM_NONE);
				@(negedge vif.pready);

			end
			$display("----------------------------------------------");
			$display("                                              ");
			$display("----------------------------------------------");
			seq_item_port.item_done();
		end
	endtask
endclass


class monitor extends uvm_monitor;
	`uvm_component_utils(monitor)

	uvm_analysis_port #(transaction) send;
    transaction tr;
	virtual apb_if vif;
  
  	covergroup apb_data;
    
    	option.per_instance = 1;
    
      	Read_Write : coverpoint tr.pwrite{
        	bins read = {0};
        	bins write = {1};
      	}

      	Addr : coverpoint tr.paddr{
        	bins valid_addr[] = {[0:31]};
        	bins invalid_addr = default;
      	}

      	Error : coverpoint tr.pslverr{
        	bins valid_trans = {0};
        	bins error = {1};
      	}
      
      	Write_Data : coverpoint tr.pwdata{
        	bins low = {[0 : 32'h3fff_ffff]};
        	bins mid1 = {[32'h4000_0000 : 32'h7fff_ffff]};
        	bins mid2 = {[32'h8000_0000 : 32'hbfff_ffff]};
        	bins high = {[32'hC000_0000 : 32'hffff_ffff]};
      	}
      
      	Read_Data : coverpoint tr.prdata{
        	bins low = {[0 : 32'h3fff_ffff]};
        	bins mid1 = {[32'h4000_0000 : 32'h7fff_ffff]};
        	bins mid2 = {[32'h8000_0000 : 32'hbfff_ffff]};
        	bins high = {[32'hC000_0000 : 32'hffff_ffff]};
      	}
      
        
      
      	Addr_cvr_write : cross Read_Write, Addr{
        	ignore_bins unused = binsof(Read_Write) intersect {0}; 
      	}
      
      	Addr_cvr_read : cross Read_Write, Addr{
        	ignore_bins unused = binsof(Read_Write) intersect {1}; 
      	}
      
      	WData_cvr_write : cross Read_Write, Write_Data{
        	ignore_bins unused = binsof(Read_Write) intersect {0}; 
      	}
      
      	RData_cvr_read : cross Read_Write, Read_Data{
        	ignore_bins unused = binsof(Read_Write) intersect {1}; 
      	}
      
      	Err_cvr_write : cross Read_Write, Error{
        	ignore_bins unused_write = binsof(Read_Write) intersect {0};
        	ignore_bins no_error = binsof(Error) intersect{0};
      	}
      
      	Err_cvr_read : cross Read_Write, Error{
        	ignore_bins unused_read = binsof(Read_Write) intersect {1};
        	ignore_bins no_error = binsof(Error) intersect{0};
      	}
      
      
    endgroup
  
  
  	
	function new(input string path = "monitor", input uvm_component parent = null);
		super.new(path,parent);
      	apb_data = new();
	endfunction

	

	virtual function void build_phase(uvm_phase phase);
		super.build_phase(phase);

		tr = transaction::type_id::create("tr");
		send = new("send",this);

		if(!uvm_config_db#(virtual apb_if)::get(this,"","vif",vif))
			`uvm_error("MON","Unable to access Virtual Interface");
	endfunction
	

	virtual task run_phase(uvm_phase phase);
		forever begin

			@(posedge vif.pclk);
			if(vif.presetn == 0)
			begin
				tr.op = rst;
				`uvm_info("MON","Reset Detected",UVM_NONE);
				send.write(tr);
			end

			else if(vif.pwrite)
			begin
				@(posedge vif.pready)
				tr.op = writed;
				tr.pwdata = vif.pwdata;
				tr.paddr = vif.paddr;
				tr.pslverr = vif.pslverr;
              	tr.pwrite = vif.pwrite;
              	apb_data.sample();
				`uvm_info("MON",$sformatf("Data Write Received From Interface: Addr = %0d, WData = %0d, Slave Error = %0b",vif.paddr, vif.pwdata, vif.pslverr),UVM_NONE);
				@(negedge vif.pready);
				send.write(tr);
			end

			else if(!vif.pwrite)
			begin
				@(posedge vif.pready)
				tr.op = readd;
				tr.prdata = vif.prdata;
				tr.paddr = vif.paddr;
				tr.pslverr = vif.pslverr;
              	tr.pwrite = vif.pwrite;
              	apb_data.sample();
				`uvm_info("MON",$sformatf("Data Read Received From Interface: Addr = %0d, Rdata = %0d, Slave Error = %0b",vif.paddr, vif.prdata, vif.pslverr),UVM_NONE);
				@(negedge vif.pready);
				send.write(tr);

			end


		end
	endtask
endclass



class scoreboard extends uvm_scoreboard;
	`uvm_component_utils(scoreboard)

	logic [31:0] addr = 0;
	logic [31:0] mem [32] = '{default:0};
	logic [31:0] data_rd = 0;

	uvm_analysis_imp #(transaction, scoreboard) rcv;

	function new(string path = "sco", uvm_component parent = null);
		super.new(path,parent);
	endfunction

	virtual function void build_phase(uvm_phase phase);
		super.build_phase(phase);

		rcv = new("rcv",this);

	endfunction

	virtual function void write(input transaction tr);

		if(tr.op == rst)
		begin
			`uvm_info("SCO","Reset Detected",UVM_NONE)
			for(int i = 0; i < 32; i++) 
        		begin
          			mem[i] = 0;
        		end	
		end

		else if(tr.op == writed)
		begin
			if(tr.pslverr && (tr.paddr > 32))
				`uvm_info("SCO","Error Successfully Detected",UVM_LOW)
			else if(!tr.pslverr && (tr.paddr < 32))begin
				mem[tr.paddr] = tr.pwdata;
				`uvm_info("SCO",$sformatf("Data Written Successfully : Addr = %0d, Wdata = %0d", tr.paddr, tr.pwdata),UVM_LOW)

			end
			else
			begin
				`uvm_error("SCO","Some Error in Detecting Illegal Address")
			end
		end

		else if(tr.op == readd)
		begin
			if(tr.pslverr && (tr.paddr > 32))
				`uvm_info("SCO","Error Successfully Detected",UVM_LOW)
			else if(!tr.pslverr && (tr.paddr < 32))begin
				data_rd = mem[tr.paddr];

				`uvm_info("SCO","Data Received",UVM_LOW);
				if(data_rd == tr.prdata)
					`uvm_info("SCO",$sformatf("Data MATCHED: Addr = %0d, Rdata = %0d",tr.paddr, tr.prdata),UVM_LOW)
				else
					`uvm_error("SCO",$sformatf("Data MISMATCH: Addr = %0d, Expected = %0d, Received = %0d",tr.paddr, data_rd, tr.prdata))
			end
			else
			begin
				`uvm_error("SCO","Some Error in Detecting Illegal Address")
			end
		end
	

	endfunction
endclass


class agent extends uvm_agent;
`uvm_component_utils(agent)
 
 	apb_config cfg;

	function new(input string inst = "AGENT", uvm_component c);
		super.new(inst, c);
	endfunction

	uvm_sequencer #(transaction) seqr;
	driver drv;
	monitor mon;

	virtual function void build_phase(uvm_phase phase);
		super.build_phase(phase);

		cfg = apb_config::type_id::create("cfg");
		mon = monitor::type_id::create("mon",this);
		
		if(cfg.is_active == UVM_ACTIVE) begin
			seqr = uvm_sequencer #(transaction)::type_id::create("seqr",this);
			drv = driver::type_id::create("drv",this);
		end
	endfunction

	virtual function void connect_phase(uvm_phase phase);
		super.connect_phase(phase);

		if(cfg.is_active == UVM_ACTIVE) begin
			drv.seq_item_port.connect(seqr.seq_item_export);
		end

	endfunction
endclass


class env extends uvm_env;
	`uvm_component_utils(env)
 
 
	function new(input string inst = "ENV", uvm_component c);
		super.new(inst, c);
	endfunction

	agent a;
	scoreboard sco;

	virtual function void build_phase(uvm_phase phase);
		super.build_phase(phase);

		a = agent::type_id::create("a",this);
		sco = scoreboard::type_id::create("sco",this);
	endfunction

	virtual function void connect_phase(uvm_phase phase);
		super.connect_phase(phase);

		a.mon.send.connect(sco.rcv);
	endfunction
endclass

class test extends uvm_test;
	`uvm_component_utils(test)

	env e;
	write_data writed;
	write_err writeerr;
	read_data readd;
	read_err readerr;
	reset_dut rstdut;
	writeb_readb wrb_rdb;
	write_read wr_rd;

	function new(string path = "test", uvm_component parent = null);
		super.new(path,parent);
	endfunction

	virtual function void build_phase(uvm_phase phase);
		super.build_phase(phase);

		e = env::type_id::create("e",this);
		
		writed = write_data::type_id::create("writed");
		writeerr = write_err::type_id::create("writeerr");
		readd = read_data::type_id::create("readd");
		readerr = read_err::type_id::create("readerr");
		rstdut = reset_dut::type_id::create("rstdut");	
		wrb_rdb = writeb_readb::type_id::create("wrb_rdb");
		wr_rd = write_read::type_id::create("wr_rd");

	
	endfunction

	virtual task run_phase(uvm_phase phase);
		phase.raise_objection(this);
		writed.start(e.a.seqr);
		#20
		`uvm_info("TEST","Write Sequence Executed",UVM_NONE)

		$display("////////////////////////////////////////////////////////////////////");
		$display("");
		$display("");
		$display("");
		$display("////////////////////////////////////////////////////////////////////");
		
		readd.start(e.a.seqr);
		//#20;
		`uvm_info("TEST","Read Sequence Executed",UVM_NONE)
		
		$display("////////////////////////////////////////////////////////////////////");
		$display("");
		$display("");
		$display("");
		$display("////////////////////////////////////////////////////////////////////");

		rstdut.start(e.a.seqr);
		#20
		`uvm_info("TEST","Reset Sequence Executed",UVM_NONE)
		
		$display("////////////////////////////////////////////////////////////////////");
		$display("");
		$display("");
		$display("");
		$display("////////////////////////////////////////////////////////////////////");
		
		writeerr.start(e.a.seqr);
		#20
		`uvm_info("TEST","Write Error Sequence Executed",UVM_NONE)
		
		$display("////////////////////////////////////////////////////////////////////");
		$display("");
		$display("");
		$display("");
		$display("////////////////////////////////////////////////////////////////////");

		readerr.start(e.a.seqr);
		`uvm_info("TEST","Read Error Sequence Executed",UVM_NONE)
		
		$display("////////////////////////////////////////////////////////////////////");
		$display("");
		$display("");
		$display("");
		$display("////////////////////////////////////////////////////////////////////");	

		wrb_rdb.start(e.a.seqr);
		//#20;
		`uvm_info("TEST","Bulk Sequence Executed",UVM_NONE)
		$display("////////////////////////////////////////////////////////////////////");
		$display("");
		$display("");
		$display("");
		$display("////////////////////////////////////////////////////////////////////");

		rstdut.start(e.a.seqr);
		#20
		`uvm_info("TEST","Reset Sequence Executed",UVM_NONE)
		
		$display("////////////////////////////////////////////////////////////////////");
		$display("");
		$display("");
		$display("");
		$display("////////////////////////////////////////////////////////////////////");

		wr_rd.start(e.a.seqr);
		#20;
		`uvm_info("TEST","Read Write Sequence Executed",UVM_NONE)
		$display("////////////////////////////////////////////////////////////////////");
		$display("");
		$display("");
		$display("");
		$display("////////////////////////////////////////////////////////////////////");

		phase.drop_objection(this);
	endtask

endclass


module tb;

	apb_if vif();
	
	apb_ram dut(.presetn(vif.presetn), .pclk(vif.pclk), .psel(vif.psel), .penable(vif.penable), .pwrite(vif.pwrite), .paddr(vif.paddr), .pwdata(vif.pwdata), .prdata(vif.prdata), .pready(vif.pready), .pslverr(vif.pslverr));
  
  	bind apb_ram apb_assertions assertion_mod (vif.pclk, vif.presetn, vif.paddr, vif.pwrite, vif.pwdata, vif.penable, vif.psel, vif.prdata, vif.pslverr, vif.pready);

	initial begin
		vif.pclk <= 0;
	end

	always #5 vif.pclk = ~vif.pclk;



  initial begin

		uvm_config_db #(virtual apb_if)::set(null,"uvm_test_top.e.a*","vif",vif);
		run_test("test");
	end


  initial begin

    $dumpfile("dump.vcd");
    $dumpvars;

  end



endmodule
